// udp_bridge_core.v

// Generated using ACDS version 22.1 915

`timescale 1 ps / 1 ps
module udp_bridge_core (
		input  wire        clk_clk,       //     clk.clk
		input  wire        ethio_enable,  //   ethio.enable
		output wire [2:0]  ethio_status,  //        .status
		input  wire [31:0] ipaddr_value,  //  ipaddr.value
		output wire [1:0]  led_export,    //     led.export
		input  wire [47:0] macaddr_value, // macaddr.value
		input  wire        reset_reset_n, //   reset.reset_n
		input  wire        rmii_clk,      //    rmii.clk
		input  wire [1:0]  rmii_rxd,      //        .rxd
		input  wire        rmii_crs_dv,   //        .crs_dv
		output wire [1:0]  rmii_txd,      //        .txd
		output wire        rmii_tx_en     //        .tx_en
	);

	wire         peridot_ethio_0_m1_waitrequest;                        // mm_interconnect_0:peridot_ethio_0_m1_waitrequest -> peridot_ethio_0:avm_m1_waitrequest
	wire  [31:0] peridot_ethio_0_m1_readdata;                           // mm_interconnect_0:peridot_ethio_0_m1_readdata -> peridot_ethio_0:avm_m1_readdata
	wire  [31:0] peridot_ethio_0_m1_address;                            // peridot_ethio_0:avm_m1_address -> mm_interconnect_0:peridot_ethio_0_m1_address
	wire         peridot_ethio_0_m1_read;                               // peridot_ethio_0:avm_m1_read -> mm_interconnect_0:peridot_ethio_0_m1_read
	wire   [3:0] peridot_ethio_0_m1_byteenable;                         // peridot_ethio_0:avm_m1_byteenable -> mm_interconnect_0:peridot_ethio_0_m1_byteenable
	wire         peridot_ethio_0_m1_readdatavalid;                      // mm_interconnect_0:peridot_ethio_0_m1_readdatavalid -> peridot_ethio_0:avm_m1_readdatavalid
	wire         peridot_ethio_0_m1_write;                              // peridot_ethio_0:avm_m1_write -> mm_interconnect_0:peridot_ethio_0_m1_write
	wire  [31:0] peridot_ethio_0_m1_writedata;                          // peridot_ethio_0:avm_m1_writedata -> mm_interconnect_0:peridot_ethio_0_m1_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata; // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;  // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire         mm_interconnect_0_pio_0_s1_chipselect;                 // mm_interconnect_0:pio_0_s1_chipselect -> pio_0:chipselect
	wire  [31:0] mm_interconnect_0_pio_0_s1_readdata;                   // pio_0:readdata -> mm_interconnect_0:pio_0_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_0_s1_address;                    // mm_interconnect_0:pio_0_s1_address -> pio_0:address
	wire         mm_interconnect_0_pio_0_s1_write;                      // mm_interconnect_0:pio_0_s1_write -> pio_0:write_n
	wire  [31:0] mm_interconnect_0_pio_0_s1_writedata;                  // mm_interconnect_0:pio_0_s1_writedata -> pio_0:writedata
	wire         rst_controller_reset_out_reset;                        // rst_controller:reset_out -> [mm_interconnect_0:peridot_ethio_0_reset_reset_bridge_in_reset_reset, peridot_ethio_0:rsi_reset_reset, pio_0:reset_n, sysid_qsys_0:reset_n]

	peridot_ethio #(
		.RXFIFO_SIZE         (4096),
		.TXFIFO_SIZE         (4096),
		.FIFO_BLOCKSIZE      (64),
		.SUPPORT_SPEED_10M   (0),
		.SUPPORT_HARFDUPLEX  (0),
		.SUPPORT_PAUSEFRAME  (0),
		.MTU_SIZE            (1500),
		.ENABLE_UDP_CHECKSUM (1),
		.IGNORE_RXFCS_CHECK  (0),
		.FIXED_MAC_ADDRESS   (48'b000000000000000000000000000000000000000000000000),
		.FIXED_IP_ADDRESS    (32'b00000000000000000000000000000000),
		.FIXED_UDP_PORT      (16241),
		.FIXED_PAUSE_LESS    (0),
		.FIXED_PAUSE_VALUE   (0),
		.SUPPORT_MEMORYHOST  (1),
		.AVALONMM_FASTMODE   (0),
		.SUPPORT_STREAMFIFO  (0),
		.SRCFIFO_NUMBER      (1),
		.SINKFIFO_NUMBER     (1),
		.SRCFIFO_0_SIZE      (2048),
		.SRCFIFO_1_SIZE      (2048),
		.SRCFIFO_2_SIZE      (2048),
		.SRCFIFO_3_SIZE      (2048),
		.SINKFIFO_0_SIZE     (2048),
		.SINKFIFO_1_SIZE     (2048),
		.SINKFIFO_2_SIZE     (2048),
		.SINKFIFO_3_SIZE     (2048)
	) peridot_ethio_0 (
		.csi_clock_clk        (clk_clk),                          //   clock.clk
		.rsi_reset_reset      (rst_controller_reset_out_reset),   //   reset.reset
		.avm_m1_waitrequest   (peridot_ethio_0_m1_waitrequest),   //      m1.waitrequest
		.avm_m1_address       (peridot_ethio_0_m1_address),       //        .address
		.avm_m1_read          (peridot_ethio_0_m1_read),          //        .read
		.avm_m1_readdata      (peridot_ethio_0_m1_readdata),      //        .readdata
		.avm_m1_readdatavalid (peridot_ethio_0_m1_readdatavalid), //        .readdatavalid
		.avm_m1_write         (peridot_ethio_0_m1_write),         //        .write
		.avm_m1_writedata     (peridot_ethio_0_m1_writedata),     //        .writedata
		.avm_m1_byteenable    (peridot_ethio_0_m1_byteenable),    //        .byteenable
		.coe_enable           (ethio_enable),                     //   ethio.enable
		.coe_status           (ethio_status),                     //        .status
		.coe_macaddr          (macaddr_value),                    // macaddr.value
		.coe_ipaddr           (ipaddr_value),                     //  ipaddr.value
		.coe_rmii_clk         (rmii_clk),                         //    rmii.clk
		.coe_rmii_rxd         (rmii_rxd),                         //        .rxd
		.coe_rmii_crsdv       (rmii_crs_dv),                      //        .crs_dv
		.coe_rmii_txd         (rmii_txd),                         //        .txd
		.coe_rmii_txen        (rmii_tx_en),                       //        .tx_en
		.aso_src0_ready       (1'b0),                             // (terminated)
		.aso_src0_valid       (),                                 // (terminated)
		.aso_src0_data        (),                                 // (terminated)
		.aso_src1_ready       (1'b0),                             // (terminated)
		.aso_src1_valid       (),                                 // (terminated)
		.aso_src1_data        (),                                 // (terminated)
		.aso_src2_ready       (1'b0),                             // (terminated)
		.aso_src2_valid       (),                                 // (terminated)
		.aso_src2_data        (),                                 // (terminated)
		.aso_src3_ready       (1'b0),                             // (terminated)
		.aso_src3_valid       (),                                 // (terminated)
		.aso_src3_data        (),                                 // (terminated)
		.asi_sink0_ready      (),                                 // (terminated)
		.asi_sink0_valid      (1'b0),                             // (terminated)
		.asi_sink0_data       (8'b00000000),                      // (terminated)
		.asi_sink1_ready      (),                                 // (terminated)
		.asi_sink1_valid      (1'b0),                             // (terminated)
		.asi_sink1_data       (8'b00000000),                      // (terminated)
		.asi_sink2_ready      (),                                 // (terminated)
		.asi_sink2_valid      (1'b0),                             // (terminated)
		.asi_sink2_data       (8'b00000000),                      // (terminated)
		.asi_sink3_ready      (),                                 // (terminated)
		.asi_sink3_valid      (1'b0),                             // (terminated)
		.asi_sink3_data       (8'b00000000),                      // (terminated)
		.coe_speed10m         (1'b0),                             // (terminated)
		.coe_halfduplex       (1'b0),                             // (terminated)
		.coe_udpport          (16'b0000000000000000),             // (terminated)
		.coe_pause_less       (8'b00000000),                      // (terminated)
		.coe_pause_value      (16'b0000000000000000)              // (terminated)
	);

	udp_bridge_core_pio_0 pio_0 (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_pio_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_0_s1_readdata),   //                    .readdata
		.out_port   (led_export)                             // external_connection.export
	);

	udp_bridge_core_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_clk),                                               //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	udp_bridge_core_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                     (clk_clk),                                               //                                   clk_0_clk.clk
		.peridot_ethio_0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                        // peridot_ethio_0_reset_reset_bridge_in_reset.reset
		.peridot_ethio_0_m1_address                        (peridot_ethio_0_m1_address),                            //                          peridot_ethio_0_m1.address
		.peridot_ethio_0_m1_waitrequest                    (peridot_ethio_0_m1_waitrequest),                        //                                            .waitrequest
		.peridot_ethio_0_m1_byteenable                     (peridot_ethio_0_m1_byteenable),                         //                                            .byteenable
		.peridot_ethio_0_m1_read                           (peridot_ethio_0_m1_read),                               //                                            .read
		.peridot_ethio_0_m1_readdata                       (peridot_ethio_0_m1_readdata),                           //                                            .readdata
		.peridot_ethio_0_m1_readdatavalid                  (peridot_ethio_0_m1_readdatavalid),                      //                                            .readdatavalid
		.peridot_ethio_0_m1_write                          (peridot_ethio_0_m1_write),                              //                                            .write
		.peridot_ethio_0_m1_writedata                      (peridot_ethio_0_m1_writedata),                          //                                            .writedata
		.pio_0_s1_address                                  (mm_interconnect_0_pio_0_s1_address),                    //                                    pio_0_s1.address
		.pio_0_s1_write                                    (mm_interconnect_0_pio_0_s1_write),                      //                                            .write
		.pio_0_s1_readdata                                 (mm_interconnect_0_pio_0_s1_readdata),                   //                                            .readdata
		.pio_0_s1_writedata                                (mm_interconnect_0_pio_0_s1_writedata),                  //                                            .writedata
		.pio_0_s1_chipselect                               (mm_interconnect_0_pio_0_s1_chipselect),                 //                                            .chipselect
		.sysid_qsys_0_control_slave_address                (mm_interconnect_0_sysid_qsys_0_control_slave_address),  //                  sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata               (mm_interconnect_0_sysid_qsys_0_control_slave_readdata)  //                                            .readdata
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
